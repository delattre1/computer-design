library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

entity memoriaROM is
   generic (
          dataWidth: natural := 13;
          addrWidth: natural := 9
    );
   port (
          Endereco : in std_logic_vector (addrWidth-1 DOWNTO 0);
          Dado     : out std_logic_vector(dataWidth-1 DOWNTO 0)
    );
end entity;

architecture assincrona of memoriaROM is

  type blocoMemoria is array(0 TO 2**addrWidth - 1) of std_logic_vector(dataWidth-1 DOWNTO 0);

  function initMemory 
        return blocoMemoria is variable tmp : blocoMemoria := (others => (others => '0'));
  begin
			  -- Inicializa os endereços: Testa JMP
			--tmp(0) := "0000000000000";  -- NOP	
			--tmp(1) := "0110000000100";  -- JMP @4	
			--tmp(2) := "0110000000101";  -- JMP @5	
			--tmp(3) := "0000000000000";  -- NOP	
			--tmp(4) := "0000000000000";  -- NOP	
			--tmp(5) := "0110000000001";  -- JMP @1	
			
			-- tmp(0)  :=  "0000000000000"; -- NOP
			-- tmp(1)  :=  "0110000000100"; -- JMP @4	 -- Deve desviar para a posição 4
			-- tmp(2)  :=  "0111000001001"; -- JEQ @9	 -- Deve desviar para a posição 9
			-- tmp(3)  :=  "0000000000000"; -- NOP	 -- 
			-- tmp(4)  :=  "0000000000000"; -- NOP	 -- 
			-- tmp(5)  :=  "0100000000101"; -- LDI $5	 -- Carrega acumulador com valor 5
			-- tmp(6)  :=  "0101000000000"; -- STA @0	 -- Armazena 5 na posição 0 da memória
			-- tmp(7)  :=  "1000000000000"; -- CEQ @0	 -- A comparação deve fazer o flagIgual ser 1
			-- tmp(8)  :=  "0110000000001"; -- JMP @1	 -- Vai testar o flagIgual depois do jump
			-- tmp(9)  :=  "0000000000000"; -- NOP	 -- 
			-- tmp(10) :=  "0100000000100"; -- LDI $4	 -- Carrega acumulador com valor 4
			-- tmp(11) :=  "1000000000000"; -- CEQ @0	 -- Compara com valor 5, deve fazer o flagIgual ser 0
			-- tmp(12) :=  "0111000000011"; -- JEQ @3	 -- Não deve ocorrer o desvio
			-- tmp(13) :=  "0110000001100"; -- JMP @12 -- Fim. Deve ficar neste laço enableWriteRet <= Sinais_Controle(11);
			tmp(0)  :=  "1001000001110"; --JSR @14	Deve desviar para a posição 14
			tmp(1)  :=  "0110000000101"; --JMP @5	Deve desviar para a posição 5
			tmp(2)  :=  "0111000001001"; --JEQ @9	Deve desviar para a posição 9
			tmp(3)  :=  "0000000000000"; --NOP	
			tmp(4)  :=  "0000000000000"; --NOP	
			tmp(5)  :=  "0100000000101"; --LDI $5	Carrega acumulador com valor 5
			tmp(6)  :=  "0101000000000"; --STA @0	Armazena 5 na posição 0 da memória
			tmp(7)  :=  "1000000000000"; --CEQ @0	A comparação deve fazer o flagIgual ser 1
			tmp(8)  :=  "0110000000010"; --JMP @2	Vai testar o flagIgual depois do jump
			tmp(9)  :=  "0000000000000"; --NOP	
			tmp(10) :=  "0100000000100"; --LDI $4	Carrega acumulador com valor 4
			tmp(11) :=  "1000000000000"; --CEQ @0	Compara com valor 5, deve fazer o flagIgual ser 0
			tmp(12) :=  "0111000000011"; --JEQ @3	Não deve ocorrer o desvio
			tmp(13) :=  "0110000001101"; --JMP @13	Fim. Deve ficar neste laço
			tmp(14) :=  "0000000000000"; --NOP	
			tmp(15) :=  "1010000000000"; --RET	Retorna para a posição 1

			return tmp;
    end initMemory;

    signal memROM : blocoMemoria := initMemory;

begin
    Dado <= memROM (to_integer(unsigned(Endereco)));
end architecture;